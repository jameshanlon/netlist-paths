module include_a(
                 input  data_i,
                 output data_o
                 );

   assign data_o = data_i;

endmodule
