module single_define(
               input data_i,
               output data_o
               );

   assign data_o = `EXPR_A;

endmodule
