// test multiple independent top levels
module top_b(
             input  data_b_i,
             output data_b_o
             );

   assign data_b_o = data_b_i;

endmodule
