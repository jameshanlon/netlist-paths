module empty_module
  (
    input in,
    output out
  );
endmodule
