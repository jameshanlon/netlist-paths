// test multiple independent top levels
module top_a(
             input  data_a_i,
             output data_a_o
             );

   assign data_a_o = data_a_i;

endmodule
